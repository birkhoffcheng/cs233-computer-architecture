module logicunit_test;
    // exhaustively test your logic unit implementation by adapting mux4_tb.v
endmodule // logicunit_test
