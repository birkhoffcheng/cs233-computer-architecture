module alu1_test;
    // exhaustively test your 1-bit ALU implementation by adapting mux4_tb.v
endmodule
