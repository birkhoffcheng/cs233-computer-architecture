//implement a test bench for your 32-bit ALU
module alu32_test;
	reg [31:0] A = 0, B = 0;
	reg [2:0] control = 0;

	initial begin
		$dumpfile("alu32.vcd");
		$dumpvars(0, alu32_test);

			 A = 8; B = 4; control = `ALU_ADD; // try adding 8 and 4
		# 10 A = 2; B = 5; control = `ALU_SUB; // try subtracting 5 from 2
		// add more test cases here!

		# 10 $finish;
	end

	wire [31:0] out;
	wire overflow, zero, negative;
	alu32 a(out, overflow, zero, negative, A, B, control);

	integer myint;
	always @(out) myint = out;
	
	initial begin
		$display("\tA\t\tB\tcontrol\t\tint\t\tout\toverflow\tzero\tnegative");
		$monitor("%d\t%d\t%d\t%d\t%d\t%d\t\t%d\t%d\t(at time %t)", A, B, control, myint, out, overflow, zero, negative, $time);
	end
endmodule // alu32_test
