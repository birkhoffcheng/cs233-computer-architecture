module blackbox_test;

endmodule // blackbox_test
