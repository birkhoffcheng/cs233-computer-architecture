//Write your test bench for sc2_block here.
//Refer to sc_block_tb.v for formatting!
module sc2_test;

endmodule // sc2_test
